library verilog;
use verilog.vl_types.all;
entity Lab6Block_vlg_vec_tst is
end Lab6Block_vlg_vec_tst;
