library verilog;
use verilog.vl_types.all;
entity P3_vlg_vec_tst is
end P3_vlg_vec_tst;
