library verilog;
use verilog.vl_types.all;
entity Arjen_Arumalingam_Lab6_vlg_vec_tst is
end Arjen_Arumalingam_Lab6_vlg_vec_tst;
